library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity Imemory is
    Port ( address : in   STD_LOGIC_VECTOR (11 downto 0);
           instruction : out  STD_LOGIC_VECTOR (31 downto 0));
end Imemory;
architecture Behavioral of Imemory is
type memory_type is array (0 to (2**12)-1) of std_logic_vector (31 downto 0);
constant memory : memory_type  := ("00101100000000000000000000001110",
"00110000000000000000000001111100",
"00100000000000000000000001000101",
"00110000000000000000000010011101",
"00100000000000000000000001000101",
"00110000000000000000000010011101",
"00100000000000000000000001000101",
"00110000000000000000000010011101",
"00100000000000000000000001000101",
"00110000000000000000000010011101",
"00100000000000000000000001000101",
"00110000000000000000000010011101",
"00100000000000000000000001000101",
"00110000000000000000000010011101",
"00110000000000000000000000010000",
"00101100000000000000000000001110",
"01010011110000000000000000000000",
"00001001111011111000011111111111",
"01001001111000000000000000000000",
"01011100000000000000000000000000",
"01011100000000000000000000000000",
"01011100000000000000000000000000",
"00100000000000110000000000001111",
"01000000000011100000000000000000",
"00001001110011100000000000001111",
"00010100011011101111111111111001",
"01011100000000000000000000000000",
"01011100000000000000000000000000",
"01011100000000000000000000000000",
"01000000000011100000000000000000",
"00000001110000110111000000000100",
"00001100011011011111111111110111",
"00110000000000000000000001101010",
"01000000000011100000000000000000",
"01000000000011100000000000000000",
"00000001110000110111000000000100",
"00001100011011011111111111110010",
"00100000000011110111000000000000",
"01001001111000000000000000000000",
"01011100000000000000000000000000",
"01011100000000000000000000000000",
"01011100000000000000000000000000",
"01000000000011100000000000000000",
"00000001110000110111000000000100",
"00010100011011110000000000011000",
"00100000000011110110100000000000",
"01001001111000000000000000000000",
"01011100000000000000000000000000",
"01011100000000000000000000000000",
"01011100000000000000000000000000",
"01000000000011100000000000000000",
"00000001110000110111000000000100",
"00010100011011110000000000010010",
"00100000000011110101100000000000",
"01001001111000000000000000000000",
"01011100000000000000000000000000",
"01011100000000000000000000000000",
"01011100000000000000000000000000",
"01000000000011100000000000000000",
"00000001110000110111000000000100",
"00010100011011110000000000001100",
"00100000000011110011100000000000",
"01001001111000000000000000000000",
"01011100000000000000000000000000",
"01011100000000000000000000000000",
"01011100000000000000000000000000",
"01000000000011100000000000000000",
"00000001110000110111000000000100",
"00010100011011110000000000000110",
"00100000000101000000000000000000",
"00101100000000000000000001001100",
"00100000000101000000000000000100",
"00101100000000000000000001001100",
"00100000000101000000000000001000",
"00101100000000000000000001001100",
"00100000000101000000000000001100",
"01010001110000000000000000000000",
"00001001110011100000000000001000",
"00100000000101010000000000001000",
"00010110101011110000000000000011",
"00000110100101000000000000000000",
"01001100000011100000000000000000",
"00101100000000000000000001100101",
"01001100000011100000000000000000",
"01010001110000000000000000000000",
"00001001110011100000000000000100",
"00100000000101010000000000000100",
"00010110101011110000000000000011",
"00000110100101000000000000000001",
"01001100000011100000000000000000",
"00101100000000000000000001100101",
"01001100000011100000000000000000",
"01010001110000000000000000000000",
"00001001110011100000000000000010",
"00100000000101010000000000000010",
"00010110101011110000000000000011",
"00000110100101000000000000000010",
"01001100000011100000000000000000",
"00101100000000000000000001100101",
"01001100000011100000000000000000",
"00000110100101000000000000000011",
"01010011110000000000000000000000",
"00011101110000000000000000000000",
"00110000000000000000000010011101",
"01001100000111100000000000000000",
"00111011110000000000000000000000",
"01010011110000000000000000000000",
"00100000000111110000000010100000",
"00110000000000000000000001111000",
"00000011111000001111100000001111",
"00110100000000000000000001101100",
"01001100000111100000000000000000",
"00111011110000000000000000000000",
"01010011110000000000000000000000",
"00100000000111010000000001100100",
"00110000000000000000000001111000",
"00000011101000001110100000001111",
"01011011101111010000000001110011",
"01001100000111100000000000000000",
"00111011110000000000000000000000",
"00100000000111110000010011100010",
"00000011111000001111100000001111",
"00110100000000000000000001111001",
"00111011110000000000000000000000",
"01010011110000000000000000000000",
"00001000000000000000000000000000",
"01001000000000000000000000000000",
"00110000000000000000000001110001",
"00100100000000000000000000111000",
"00110000000000000000000010010001",
"00110000000000000000000001110001",
"00001000000000000000000000000000",
"00100100000000000000000000001110",
"00110000000000000000000010010001",
"00110000000000000000000001110001",
"00001000000000000000000000000000",
"00100100000000000000000000000001",
"00110000000000000000000010010001",
"00110000000000000000000001110001",
"00001000000000000000000000000000",
"00100100000000000000000000000110",
"00110000000000000000000010010001",
"00110000000000000000000001110001",
"01001100000111100000000000000000",
"00111011110000000000000000000000",
"01010011110000000000000000000000",
"00001001111011111111100000000000",
"00001000000000000000000011111111",
"00000001111000000111100000000101",
"00100101111011110000000100000000",
"01001001111000000000000000000000",
"00110000000000000000000001110001",
"00001001111011111111111011111111",
"01001001111000000000000000000000",
"00110000000000000000000001110001",
"01001100000111100000000000000000",
"00111011110000000000000000000000",
"01010011110000000000000000000000",
"00001001111011111111100000000000",
"00001000000000000000000011111111",
"00000001111000000111100000000101",
"01001001111000000000000000000000",
"00100101111011110000010100000000",
"01001001111000000000000000000000",
"00110000000000000000000001110001",
"00001001111011111111111011111111",
"01001001111000000000000000000000",
"00110000000000000000000001110001",
"01001100000111100000000000000000",
"00111011110000000000000000000000",
"01010100000000000000000000000000", -- hlt
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"00000000000000000000000000000000",
"11111111111111111111111111111111",
"11111111111111111111111111111111",
"00000000000000000000000000000000"); --end at 4105 
-- hlt is "01010100000000000000000000000000"
begin
		instruction <= memory(to_integer(unsigned((address))));

end Behavioral;

